module elevator(clk, rst, inG, in1, in2, in3, in4, in5, in6, in7, up, down, open, close);

input clk, rst, inG, in1, in2, in3, in4, in5, in6, in7;
output up, down, open, close; 





endmodule